module vduckdb

pub fn library_name() {
	println('vduckdb')
}